parameter ADDR_TRIG_COUNT     = 0;
parameter ADDR_PULSE_COUNT    = 1;
parameter ADDR_DECIMATION     = 2;
parameter ADDR_DETECT_OFFSET  = 3;
parameter ADDR_TRIG_OFFSET    = 4;
parameter ADDR_CUR_TRIG       = 5;
parameter ADDR_AVERAGE_POWER  = 6;
parameter ADDR_ENABLE         = 7;
parameter ADDR_LOW_TRIG_TICKS = 8;
parameter ADDR_STOP           = ADDR_LOW_TRIG_TICKS;